logic [31:0] data = '0;
